`timescale 1ns / 1ps

module clz(
    input [31:0] in_data,
    output reg [5:0] zeros
    );
    always@(*)
    begin
    casex(in_data)
        32'b1???_????_????_????_????_????_????_????:zeros<=6'd0;
        32'b01??_????_????_????_????_????_????_????:zeros<=6'd1;
        32'b001?_????_????_????_????_????_????_????:zeros<=6'd2;
        32'b0001_????_????_????_????_????_????_????:zeros<=6'd3;
        32'b0000_1???_????_????_????_????_????_????:zeros<=6'd4;
        32'b0000_01??_????_????_????_????_????_????:zeros<=6'd5;
        32'b0000_001?_????_????_????_????_????_????:zeros<=6'd6;
        32'b0000_0001_????_????_????_????_????_????:zeros<=6'd7;
        32'b0000_0000_1???_????_????_????_????_????:zeros<=6'd8;
        32'b0000_0000_01??_????_????_????_????_????:zeros<=6'd9;
        32'b0000_0000_001?_????_????_????_????_????:zeros<=6'd10;
        32'b0000_0000_0001_????_????_????_????_????:zeros<=6'd11;
        32'b0000_0000_0000_1???_????_????_????_????:zeros<=6'd12;
        32'b0000_0000_0000_01??_????_????_????_????:zeros<=6'd13;
        32'b0000_0000_0000_001?_????_????_????_????:zeros<=6'd14;
        32'b0000_0000_0000_0001_????_????_????_????:zeros<=6'd15;
        32'b0000_0000_0000_0000_1???_????_????_????:zeros<=6'd16;
        32'b0000_0000_0000_0000_01??_????_????_????:zeros<=6'd17;
        32'b0000_0000_0000_0000_001?_????_????_????:zeros<=6'd18;
        32'b0000_0000_0000_0000_0001_????_????_????:zeros<=6'd19;
        32'b0000_0000_0000_0000_0000_1???_????_????:zeros<=6'd20;
        32'b0000_0000_0000_0000_0000_01??_????_????:zeros<=6'd21;
        32'b0000_0000_0000_0000_0000_001?_????_????:zeros<=6'd22;
        32'b0000_0000_0000_0000_0000_0001_????_????:zeros<=6'd23;
        32'b0000_0000_0000_0000_0000_0000_1???_????:zeros<=6'd24;
        32'b0000_0000_0000_0000_0000_0000_01??_????:zeros<=6'd25;
        32'b0000_0000_0000_0000_0000_0000_001?_????:zeros<=6'd26;
        32'b0000_0000_0000_0000_0000_0000_0001_????:zeros<=6'd27;
        32'b0000_0000_0000_0000_0000_0000_0000_1???:zeros<=6'd28;
        32'b0000_0000_0000_0000_0000_0000_0000_01??:zeros<=6'd29;
        32'b0000_0000_0000_0000_0000_0000_0000_001?:zeros<=6'd30;
        32'b0000_0000_0000_0000_0000_0000_0000_0001:zeros<=6'd31;
        32'b0000_0000_0000_0000_0000_0000_0000_0000:zeros<=6'd32;
     
        endcase
    end
endmodule
